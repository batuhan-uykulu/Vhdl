library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity alextender is
--  Port ( );
end alextender;

architecture Behavioral of alextender is

begin


end Behavioral;
